localparam MAX_BITS = 256;
localparam MAX_BITS_LOG2 = 8;
localparam LOOPBACK_QUEUE_COUNTER_LEN_LOG2 = 20;
localparam LOOPBACK_QUEUE_LEN_LOG2 = 10;
localparam LOOPBACK_MESSAGE_LEN = 32;
localparam CHIP_ID_LEN = 16;
localparam SFO_CTR_LEN = 1024;
localparam SFO_CTR_LEN_LOG2 = 10;
localparam SFO_CTR_INCR = 1;
localparam JITTER_INCR = 10;
localparam JITTER_MIN = 100;
localparam MAX_CHIPS_PER_SYMBOL_LOG2 = 6;
localparam CORR_WAIT_LEN_LOG2 = 15;
localparam ASSIGNMENT_SKIRT_WIDTH = 30;
localparam SKIRT_WIDTH = 2;
localparam SKIRT_WIDTH_LOG2 = 1;
localparam RECHARGE_CYCLES = 85;
localparam SYMBOL_CYCLES = 4;
localparam ESAMP_WIDTH = 20;
localparam GLOBAL_SEARCH_LEN = 3;
localparam GLOBAL_SEARCH_LEN_LOG2 = 2;
localparam PULSE_SEPARATION_LOG2 = 1;
localparam PRIMARY_FFT_LEN = 1024;
localparam PRIMARY_FFT_LEN_LOG2 = 10;
localparam PRIMARY_FFT_LEN_DECIM_LOG2 = 6;
localparam PRIMARY_FFT_WIDTH = 16;
localparam PRIMARY_FFT_MAX_LEN = 1024;
localparam PRIMARY_FFT_MAX_LEN_LOG2 = 10;
localparam PRIMARY_FFT_MAX_LEN_LOG2_LOG2 = 4;
localparam PRIMARY_FFT_DECIM_LOG2 = 4;
localparam PRIMARY_FFT_DECIM = 16;
localparam PRIMARY_FFT_MAX_LEN_DECIM_LOG2 = 6;
localparam PRIMARY_FFT_MAX_LEN_DECIM_LOG2_LOG2 = 3;
localparam SEARCH_COUNTER_LEN_LOG2 = 3;
localparam SECONDARY_FFT_LEN = 2048;
localparam SECONDARY_FFT_LEN_LOG2 = 11;
localparam SECONDARY_FFT_MAX_LEN_LOG2 = 11;
localparam SECONDARY_FFT_MAX_LEN_LOG2_LOG2 = 4;
localparam FFT_HIST_LEN = 2097152;
localparam FFT_HIST_LEN_LOG2 = 21;
localparam FFT_HIST_LEN_DECIM = 131072;
localparam FFT_HIST_LEN_DECIM_LOG2 = 17;
localparam NUM_CORRELATORS = 16;
localparam NUM_CORRELATORS_LOG2 = 4;
localparam NUM_METADATA = 7;
localparam NUM_METADATA_LOG2 = 3;
localparam OVERSAMPLING_RATIO = 16;
localparam OVERSAMPLING_RATIO_LOG2 = 4;
localparam NUM_DECODE_PATHWAYS = 5;
localparam NUM_DECODE_PATHWAYS_LOG2 = 3;
localparam PN_SEQ_LEN = 15;
localparam PN_SEQ_LEN_LOG2 = 4;
localparam SFO_INT_WIDTH = 16;
localparam SFO_FRAC_WIDTH = 16;
localparam SFO_FRAC_RANGE = 65536;
localparam SFO_SEQ_LEN_LOG2 = 7;
localparam SFO_SEQ_LEN = 72;
localparam NUM_HARMONICS = 45;
localparam NUM_HARMONICS_LOG2 = 6;
localparam RESAMPLE_INT_WIDTH = 16;
localparam RESAMPLE_FRAC_WIDTH = 15;
localparam CORR_WIDTH = 32;
localparam CORR_EXPONENT_WIDTH = 6;
localparam CORR_MANTISSA_WIDTH = 26;
localparam CORR_METADATA_WIDTH = 64;
localparam FFT_SHIFT_WIDTH = 6;
localparam [255:0] SFO_INTS = {16'd22,16'd22,16'd22,16'd22,16'd22,16'd22,16'd22,16'd22,16'd22,16'd22,16'd22,16'd22,16'd22,16'd22,16'd22,16'd22};
localparam [255:0] SFO_FRACS = {16'd22875,16'd22163,16'd21450,16'd20738,16'd20025,16'd19313,16'd18600,16'd17887,16'd17175,16'd16462,16'd15750,16'd15037,16'd14325,16'd13612,16'd12900,16'd12187};
localparam [255:0] N1S = {16'd4,16'd4,16'd4,16'd4,16'd4,16'd4,16'd4,16'd4,16'd4,16'd4,16'd4,16'd4,16'd4,16'd4,16'd4,16'd4};
localparam [239:0] N2S = {15'd3883,15'd3949,15'd4014,15'd4080,15'd4146,15'd4212,15'd4278,15'd4344,15'd4410,15'd4477,15'd4543,15'd4609,15'd4676,15'd4742,15'd4808,15'd4875};
