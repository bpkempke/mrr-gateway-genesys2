localparam GIT_VERSION=28'h404c26d;
